`include "AXI_define.svh"

module Arbiter_A()

endmodule
