`include "AXI_define.svh"
module Default_Slave(
	HandShake.in HSAR_SD,HandShake.in HSAW_SD,HandShake.in HSW_SD,
	HandShake.out HSR_SD,HandShake.out HSB_SD,
	output [1:0]logic RRESP_SD,output [1:0]logic BRESP_SD
)



endmodule
