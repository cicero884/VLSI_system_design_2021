`include "AXI_define.svh"
module Default_Master(
	//AR
	HandShake.out AR,HandShake.out AW
	//R
	//AW
	//W
	//B
);

endmodule
