`ifndef CPU_DEFINE_SVH
	`define CPU_SVH
	
	`define CPU_ADDR_BITS 14

	`define sig_Rs2 24:20
	`define sig_Rs1 19:15
	`define sig_Funct3 14:12
	`define sig_Rd 11:7
	`define sig_Opcode 6:0

`endif
